���Z     @  I   I�      Y  &                                       
    J                                                    !   �   �� 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access  �                   .       ,       )       H       �       W#       `:       �-     "�     #L     $B     +�     C�     D     E�     FZ     H#     I)     J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �0    !� BuildAll!� 0!� IDH_Contents!� Copyright � by AlexCo@     	  � 1001   �  ��:[     �  �� Et     �	 ��������"   �   ���� 
`  , 3 L     � Topic@IDH_Index  �    �I   ), , , (192,192,192), 0!�3 "Index", ( 511, 0, 511, 1023), ,$   511), , , (192,192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023%   0, 1023, 511), , , (192,192,192), 0!�. "", ( 0, 511, 1023, &    "", ( 64, 64, 832, 832), , , (192,192,192), 0!�, "", ( 0, '   6 "���������� ����������� ����", , , , (192,192,192), 0!�-(   �  _� 	   -          � F1ProjectWindowsf-�  O !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�    �, ����������� �����,(Global), 0,<IDH_Schemes>!�  !�      -   n   �� 	   .          � F1ProjectGlossary> -�   !J   �  !� 0!� 0!� No!�  !� ���������� ����������� ����!� /   rp. 1998!�  !�  !� f:\work\diplom\res\diplom.ico!� 0!�  !6    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              A   Params /Link /Macro /Play /popup/Text ���������� ��������� 2   Play /popup/Text �������� ������ ������L�L, /Jump IDH_Calc3   ��������� ��������L�L, /Jump IDH_BrigEditor /Link /Macro /4   nk /Macro /Play /popup/Text ����� ���������� ��������� ����    ere  
� �                                                6   t ������� ����!�, /P /Just L /Text Insert Menus help text h7   ������ T�     �  �� 	d�   Y -�   !� /T N /Just M /Tex8     	  � 1004   �  ��:[     �  �� Ew     � ������� �  (  ��� 
�  . 5 N     � Topic@IDH_HotKeys  �   �   ��� ����� ������������ �������� ������������/�������������;   ������ ������� �����������������.��������� �� ������������.<   �������� ����� �����������. ����� ������� ������� � �������=   � ������� � ����� �������� ����� � ������������ ��� �������   ��������!� /Z N /Style /Just L!� /X /Style /Just L  
} ?   ��� T�     �  �� 	d�   R -�   !� /T N /Just M /Text ��   ���������� ��������L�L, /Jump IDH_SimplifyMode /Link /MacroQ    !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -B   ial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None ,C   0 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , ArD   ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  12E   ,  0 , Shade , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 F    Title , Courier ,  18 ,  120 ,  250 ,  40 ,  40 ,  1 , -1 G   ?'  *� 	   ,          � F1ProjectStyle2'-�  � !�I   , (192,192,192), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�      1!�  !�  !�  !�                                            L   )�B�B,/Link /Macro /Play /Popup/Text �������� ���������� � M   ������� �������L�L, /Jump IDH_EditorSchemes /Link /Macro /PN   lay /popup/Text �������� ����������� ����L�L, /Jump IDH_EO   ditOfSchema /Link /Macro /Play /popup/Text ����� ����������P   ���� ������L�L,/Jump /Link /Macro /Play /Popup/Text �������5    ����������� ������������� ������L�L, /Jump IDH_AssPCs /LiB`   1 ,  0 , None , !�K Paragraph , System ,  10 ,  180 ,  250 a   ading , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -R     180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub HeS    20 ,  0 , -1 ,  0 , None , !�L Sub Heading , Arial ,  12 ,T   0 , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 , U   ading , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  V   12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H HeW   ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  X   , -1 , -1 , None , !�H Heading , Arial ,  12 ,  180 ,  250 Y   ading , MS Sans Serif ,  12 ,  180 ,  250 ,  60 ,  20 ,  1 Z   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�P He[    20 ,  60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  \    ,  0 , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 , ]   Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0^     10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J _   ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,Np   1 , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  4q     0 , None , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 b   paced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,c     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Sd   0 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,e    , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  6f   rial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , Noneg   250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Ah    ,  0 ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  i   �L Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10j    ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !k   ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Ariall    , -1 , None , !�M Jump Label , System ,  10 ,  180 ,  250 m   b Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1n   12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Suo   0 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  B�   ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Couri�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�T Bitmap Jump Lar    ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 , s   Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0t    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap u    0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 , v   Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 , w    24 ,  180 ,  250 ,  20 ,  60 ,  1 , -1 ,  0 , Shade , !�Q x   0 ,  0 ,  0 ,  0 , None , !�T Bitmap Paragraph , Courier , y   , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  6z   note , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 {    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Foot|    20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8}    0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 , ~   !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,    er ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,    bel , System ,  10 ,  180 ,  250 ,  20 ,  60 ,  10 ,  0 ,  �   one , !�R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  �   ns Serif ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , N�   ,  60 ,  0 ,  0 ,  0 , None , !�Z Enumerated Bullet , MS Sa�   ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20 �   G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Arial�    ,  0 ,  0 ,  0 , None , !�G Bullet , Arial ,  10 ,  180 , �    !�O Bullet , MS Sans Serif ,  10 ,  250 ,  250 ,  20 ,  60�   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,�   20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Ar�   one , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  �    , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , N�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label�   0 , None , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  25�   20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Ar�   ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M�    10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial �    0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 , �    Leaf , System ,  12 ,  440 ,  250 ,  10 ,  10 ,  1 ,  0 , �    180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�N Outline�   0 ,  0 ,  0 ,  0 , None , !�M Outline Node , Arial ,  10 , �   e , !�M Outline Node , Arial ,  10 ,  180 ,  250 ,  10 ,  1�    Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�    250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Node ,�   ,  0 ,  0 , None , !�M Outline Node , Arial ,  10 ,  180 , �   Outline Node , System ,  12 ,  180 ,  250 ,  10 ,  10 ,  0 �     10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N �    60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,�    !�R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 , �   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,��    Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 �   ter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1�   80 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Let�    -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,  1�   Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 ,�     180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index �   0 , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,�   ex Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  �   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�S Ind�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  1�   ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  25�    , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�     10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E �    250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,�   ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  440 , 6�    ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 �   60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  18�   , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  �   bel , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 �    ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter La�   one , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250�    , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , N�    20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter Label�    , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250 , �   Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None�    ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary Letter Label , �   0 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20�    !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  �   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,�   0 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Ar�   ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  18�   0 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary ,�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , �   ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,�     0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 �    , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�    Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial �   0 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 , �   0 , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  6�   Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �     10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F �   250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,�    0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 ,  �   e , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 , �    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�    , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1�   �;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None�   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�     0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,�   e , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 �    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table ,�   20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 , �     0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 ,  �    , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 , �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  �    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  �    ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  , �   , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1 �   ;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None �     , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �    0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 , �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 �    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0B   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,�   ��������L�L, /Jump IDH_Schemes /Link /Macro /Play /popup/Te�   xt ����������� ����� ������L�L, /Jump IDH_PE /Link /Macro  p/Text �������� ���� ��������� ����L�L,/Jump /Link /Macro �   up/Text ����������� �����L�L,/Jump /Link /Macro /Play /Popu�   k /Macro /Play /Popup/Text �����B�B,/Link /Macro /Play /Pop�   L,/Jump /Link /Macro /Play /Popup/Text ������L�L,/Jump /Lin�   �����������L�L,/Jump /Link /Macro /Play /Popup/Text ���L��   opup/Text ����L�L,/Jump /Link /Macro /Play /Popup/Text ����   ay /Popup/Text ������� �����L�L,/Jump /Link /Macro /Play /P�    /Play /popup/Text ����� ������ ������B�B,/Link /Macro /PlK    /Play /popup/Text ����� ��������������� (�������� ��������    �                                                          9   �   ��� 
W  , 3 L     � Topic@IDH_Menus  �    �#   0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 , 6�   /Link /Macro /Play /popup/Text ����������� ���������� �����   �����B�B,/Link /Macro /Play /Popup/Text �������������� ����   /Macro /Play /Popup/Text ��������� ������ ������ ������ �  �������� ������ ������ �������������� ������L�L,/Jump /Link  t ������� �������L�L,/Jump /Link /Macro /Play /Popup/Text �  �� �������� ��������L�L,/Jump /Link /Macro /Play /Popup/Tex�  :\work\diplom\doc\s_hot.wmf /Macro /Play /Popup /Just L  
	  	  ��� 
E / 6 O     � Topic@IDH_Contents  �  
    �  	  � 1000   �  ��=^     �  �� Hx     �
 �����  ������� W�     �  �� 	g	  ~-�   !�B /R N /Link f:\wo  rk\diplom\res\btm_app.bmp /Just M /Text ����������!�./O /J  ust L /Cols 1 /Rows 29 /Type O /Text B�B,/Link /Macro /Play   /Popup/Text ����� ���������L�L, /Jump IDH_Needing /Link /M  acro /Play /popup/Text ����������L�L, /Jump IDH_Interface    ��������� ��������B�B,/Link /Macro /Play /Popup/Text ����  /Play /Popup/Text ���� ��������� ���� ��� ������ ����������6$  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   ������ �����������, � ����������� - �������� � ������ � ���    Play /popup/Text ������  
� �                           X  �* /H /Just L /Text ���������� ���� ���������!�� /P /Just L  ����� �������� ����� ���� "���" ��� ��������� ������ ����.!  ����. ��������� ����������� ��������� ���� � ��������. ����   ����� ������� � ����� ������������� �����;!�� /B /Just L /  Text ����������� ���������� ���� ����� �� ����� �����������   ��� ����������� ����� ������ � �������������� ����������� <  ���������� ��������� �����;!�M /B /Just L /Text �������� ��   �������� MDI-���� ������������ ������ � �������� ���������  acro /Play /Popup /Just C!�
 /N /Just L!�� /P /Just L /Text  ����� ����, ������ � ������� �������������. �������������� B  ���������� ����� ��������� ����������:!�] /L /Jump IDH_Edit  ������ �������� ��������L�L, /Jump IDH_Index /Link /Macro /  ���L�L, /Jump IDH_HotKeys /Link /Macro /Play /popup/Text �0    �  	  � 3012   �  ��?`     �  �� J�     � ���  �����:!�\ /B /Just L /Text ���������� �������� �����������    0 ,  0 ,  0 ,  , !�                                        �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�4  ������� ��������� ������ ����� ��������� ��� �������  . ���%  � �����  .  ���� ����� �������� �� ����������, �� ����� ���&   ������ ���������.������� ��������� ������ ������� ��������'  � ����� ��������� ������. ������ �������� ��� ������ � ����!    {��� 
J 1 8 Q     � Topic@IDH_BrigEditor  �  .  N /Just M /Text ����� ������ �����!��/P /Just L /Text ���*  ���� ������ ������� [�     �  �� 	k�  �-�   !�& /T +      �  	  � 3011   �  ��Ab     �  �� L�     � �,  �  ���� 
" 3 : S     � Topic@IDH_SimplifyMode  �(  ���� � ���� ����� ������������ ����� ���� �����.������, ���"   N /Just M /Text �������� ������ ������!�� /P /Just L /Text/  ����� ������ �������� Y�     �  �� 	i	  h-�   !�) /T"  �������� ��������������.����������  ��������� ������� � ���A  �� ��� ������� � ��������� ���������� ���������� ���������.2  �������� ��������� ������������� ������������� ������������3  ����������� ����� �� �����;!�� /B /Just L /Text ��������� 4  ����� �������� ���������� ��������������� �������� ������ 5  ����� ������� ������ ���� ��� �������;!�h /B /Just L /Text 6  ��� � ������������������� ��������� � ����������� ��� �����7  ����� ���������;!�� /B /Just L /Text ����� ����������� ����8  ���������� ��������� ���� � ��������� ����������� ��������9   �� ���������� ����;!�n /B /Just L /Text ����� �������� ���:  st L /Text ������������ ����������� ����������� �����������;  �������� ����������� ��������� ����������� ����;!�U /B /Ju>  ����� ������� ��������������� ������������ ����������������?  � ������ �� ��������� ������� �������� ������������� ������@  ��� � ��������� �������. ������������ �� ������ ���������� 1  ���������. ������ ������������ ��� ������������� � �������K  !�H /P /Just L /Text � ���������� ������ ��� ����� ��� ����Q  orSchemes /Link /Macro /Play /popup /Just L /Text �������� D  ���������� ����� ���������������� ���������. �������� �����E  ��� ����������� �����, ������������� ������� � �����������  ���� ������.!�D /I /Jump /Link f:\work\diplom\doc\s1.wmf /M    �                                                         F  �2 /E /Just L /Text ����� ��������� �� ����� � �����.  
� G  ����� �������;!�( /E /Just L /Text ����������� ����������;!H  � ������� ������� � �����;!�+ /E /Just L /Text ��������� ��I  ������� � 1/���;!�A /E /Just L /Text �������������� �������J  ���� �����������:!�6 /E /Just L /Text ������������� ������ M  _  ��� 
$ . 5 N     � Topic@IDH_Needing  �   N   �  	  � 1005   �  ��<]     �  �� Gw     �
 ������O  ������ V�     �  �� 	fV  �-�   !� /T N /Just M /TexP  t ����������!��/P /Just L /Text ����� ���������� �������� =  ������������ ��� ������ ����������� ������������� ���������_  ����������� ����!�V /L /Jump IDH_BrigEditor /Link /Macro /a  ����� ������ �������� �������: ���� ���.��������� ������ �R  ����� �������� �������;!�k /B /Just L /Text ��������� ����S  t ��������� ���������� ������ �������� �������: ���� ���.�T  ���� �������: ���� ���.������ �������;!�b /B /Just L /TexU  ����� ������� �����������:!�E /B /Just L /Text ��������� ��V  �����, ��� ��� �� ������������ � �������� MDI-����. ��� ���W   /Text ������� ��������� ���� ������������ �� ������ �������    �  	  � 1002   �  ��>_     �  �� I�     � ����[  �  
��� 
H 0 7 P     � Topic@IDH_Interface  �  \    �  	  � 1002   �  ��>_     �  �� I�     � ����`  ������� ������������ X�     �  �� 	h�  �-�   !�) /T     ������� ������� ����������� �����  
� �                 ]  p IDH_SimplifyMode /Link /Macro /Play /popup /Just L /Text ^  Play /popup /Just L /Text �������� ������ ������!�d /L /JumC  N /Just M /Text ����������� ����������!�� /P /Just L /Text p  ������� �������;!�l /B /Just L /Text ��������� �������� ��c  ��� ������ � �����-����� ����������. � ��������� ������ ���d  ������ ���������� ����������� ������ ����� ������� �����. �e  ���� ���������� �� ����� ��������.!�F /I /Jump /Link f:\worf  k\diplom\doc\hint.wmf /Macro /Play /Popup /Just C!�) /H /Jug  st L /Text ������ ����������� �����!�u/P /Just L /Text ���h  ���� ��� ������ ��������� �����: ������ � �����������. ��� i  ������������� ����� ���� ���.����������� ��������. � ������   ������ ���������� ������������ ���������������� � ��������y  ��� ������!�/ /B /Just L /Text ������� ����� �������� Ctrl+j  ������, �����.����� ����������;!� /H /Just L /Text ����k  ������� ������������ � ����� ����������: ���� �����.������l  ����� �������: ���� �����.�������;!�p /B /Just L /Text ��m  �: ���� �����.�����;!�E /B /Just L /Text ��������� ������n  �� ������;!�B /B /Just L /Text ��������� ������������ ����o  ������� ������ �������� �������: ���� ���.�������� �������b  ����������� ����������� ������������� ������� ���� � ������  ���� �������� ���������� - ��������� �������� ������� �����r  � ����� ������ �����-���������);!�y /B /Just L /Text ��� ��s   (��� �� ����� ������ � ��������� ������ �� ����� ������� �t   �����. ������ �������� ��� ����-���������� ��������� ������  ��� ����� ���� �����.��������.!�^ /B /Just L /Text ������v  Text �������� (���� ��� ��������) ������ ����������� ������w   ������ ����� ���� ����.��������� ������.!�g /B /Just L /x  N.!�` /B /Just L /Text  ���������� (���� ����) ������ �����{  ext ����������� ����� ������� �� ������������ ������������|  ��. ������� ��� ������ ����� ���� � �� ������ ������ �� ���}  ��� ������������. ������� ������ �������� ���������� 1.1. �~  �� ����������� ���������� ����������� �������� ����� � ����  �� ���������� � 1.1. ��� ����������� �������� ������ �������  �������� �� ��������� �������������� �������� - ���������� q  � ������ ������� ������ ���������������� ��� ��������. ��� ��   ��� ��������� ������������ ����������;!�� /B /Just L /Text�  ��� �����-���� ����� � ����� ������� � ����� ������. ����� �  ������������� ���������� ������������ ������������ ���������  ������������ � ����� (����������� � ������ ����������). ����  ���, ���� � ���� ���� �� ������ ������ �� ���������. и��� �  � �������� � ���� ����� ������� �����.������� �������� �����  ��� ������� � �� ���������� ����-����� ���������� ���������  ���� � ��������� �����. ����� ������� ����� ���� ��������� �  � ����� ������ �����-���������. ������ ���������� ����������  �������� ���� � ��� ������ ��� ������ ��� ��������� ����� ��  ������.!��/P /Just L /Text ����-���������� �������� �������  ��� ��������� ������-���� ����� ����� ������ ���� ����������  ����. ��-������, ���� ����-���������� ��������������, �� � �   ���������� �������������� ���������������� � �� ������ ���z   - �������� ����� ���� �����.������������.!�}/P /Just L /Tu  �� ����� ���� ����� (����-���������� 1.1) � �� ����� �������G    �  	  � 1000   �  ��=^     �  �� Hx     �
 ������  ust L /Text ����������!�� /P /Just L /Text ������������ ����  ����� � �������������� ����. ������ ����� ������� �������� �  ������ � ������ �������������� �����. ���� ����� �������, ��  ���� ������ ��������, �� ������� ������ ����� � ������ "����  ����" ���������� ������ ����������.!� /H /Just L /Text ����  ��� �����!�0/P /Just L /Text �������������� � �������������  � ����������� ������������. ������ ����� ������ ������� ���  ��� ������� ���� ����.��������� ������. �� ����� �����������  �� ������������ ����� (�����.�����). ��� ������������ �����>   ��� ����� ������������ ������������� ���������. ��� �������    � �                                                       �   �  	  � 1003   �  ��<]     �  �� G�     � �������  � �������� ��������� V�     �  �� 	f   -�   !�* /T   N /Just M /Text ������� ������� �������!�G /I /Jump /Link fH    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   !�- /T N /Just M /Text �������� ����������� ����!� /H /J�   ��� ���� ����������� �����.!�� /B /Just L /Text ����������  ��� � ������� ����� ����������� ���� "��������".!��/B /�  �������� ����� ������������� ����� ���� �����.��������� ���  ��. � ���� ������ ��� ���� ���������.!�� /B /Just L /Text ��  ��-����� ���������� �������� ���������� �����, ��� ����� ���  ����� ������������ �������� � ����� ����� ���������� ��� ���  �������� ����� ����� ����-����� ����������. ��� ���������� �  ���������� ���������. ��� ������� ���� ����� ������������ ��  ���������� �������� � ����� � ��������� �� ����� � ������ ��  /B /Just L /Text ��������� ���������� ������������ ������ ��  ���.������������ ���������� ���������� ������ �������.!���  ���� ������.!�b /B /Just L /Text ��������� ����� � ���� ���  ���� ����� � ������ ��������� ��������� ����� ��������� �� �  �    �  	  � 3008   �  ��Bc     �  �� M�     � �  �������� ����������� ������ \�     �  �� 	la  �-�  !�  ��.�������� �������� ����� ������� ���� ����� Clipboard.�  ����� ���� ��������� ����� ����� ����.��������� �������� ��  ��.������ ����� ���������� � ������������ �����. ����������  �������� �������.!��/B /Just L /Text ����� ����� ���� ����  �������� ���������������, �� ���� ������� � ��������� ������  !�� /B /Just L /Text ���� ��������� ��������� ������ � �����   ��������� �� ������ ��������� ������� ����� � �����������.�  �����.�� � ������� �����.��������� �����. ��� ����������  ��. ����� �������� ��� ����� ����� ���� ��������������.����  ������� ��������� ������ ��� ������� ���������� ������� ����  ��� ���� ��� ��������). ��������� ���������� ���������� ����  ��� ����� ����������� ���� "��������" (������� ������ ����  Just L /Text ��������� ����������� �������������� ���������  ���� ������ ������� �� ��������� (������ �������).!�� /B /�  Just L /Text ����������� � �������. ����� ���� ����������  �����.����������, ��������������.��������, �������������  ����. �� �����.������ ������� ������� � ����� ������ ��  �� ������������ ������������. ��� ����� ���� �������� ������  �).!�Z/B /Just L /Text ������������ ��������� �����. ����  �������� ������������ ������ ��� ������ ��������� (�� ������  ������. ��������� ��������������� ���������� �������� �����  ������ �����. �������� ����� ���� ��������������.��������     /Play /popup /Just L /Text �������������� �����.  
� �  �  xt ������ �����;!�W /K /Jump IDH_EditOfSchema /Link /Macro�  Jump IDH_SimplifyMode /Link /Macro /Play /popup /Just L /Te�   /Text ���������� ��������� ������������� ��������;!�P /K /�  �:!�h /K /Jump IDH_AssPCs /Link /Macro /Play /popup /Just L�   ���� "�����".!�) /H /Just L /Text ����� ��� ������ ������  �� ���� �����. ��� ���� ����� ������� ����� ����� ����������  �� �����. ����������� ����� ���� �������������, ������������  ����� ������ ��������� ������ ����� ��������� �������� �����  ���� ������� ��� ������ ������ ��������� � ������� ������. 6�  � ���� � ����� ������� � ����� �� ������ ����� �������, ����   ����� ��������� ������ �������� �������. ��� ������ ���� ��  �� ���� "��������", � ����������� ���������� ��� ���������  ���������� ��� ������� ����������. �������� ����� ����������  �������� ��������� ������������ ���������� � ������������ ��  ����.!��/B /Just L /Text ��������� ������� ���������. �  ������� ������� �����.��������� �����, �����.��������� ��  ������������. ��� ��������� ��������� ���������� �������� �  �������� � �������.!�� /B /Just L /Text ��������� Z-�������  "���������"). ��������� ������������ ��� � ������������� �  ��� ����� ����� ��������� ������ �������  � ��������� ���� �  � �����) � ����������� ������� �����.������������ (������   ������������� ����� ������������ ����� (�����.������������   �����.��������� �� ������������. ��� ������� ������������  , ������� ������������ � ������� ����� ��������������� �����  �� ����� ������ ���� ���������� ������������ � �����. ������  ������ ��� ������ ���������� �������� ��������� ��� ��������  ���� ����� ���� ������ �� ���������� ��������� ��� �� �����  �����. �������� ����� ���� ��������������.�������, ������  ���������.������� ��, ����� ������ � �������� DEL - ����  j  uk�� 
C 4 ; T     � Topic@IDH_EditorSchemes  �  ��� ���� �� ������ �� ����);!�� /B /Just L /Text ����� ����    �������� ����� � �������� ��� ��������������.  
� �      �  ��� "�����". ����� ����������� ��� ������ ���������� ����  ����� ������ ��� ��������. ����������� ����� ����������� ��  ��������� ������ �������� �������.!�� /B /Just L /Text ����  ��������� ��������, �����. ��������� �������� ������ ����� �  ��� �������: ����������� ��������������, ��������� �����, �  � ������� ��� ������ ��������. ����� �������� ������ �������  ���. ��� ��������� ������� ������� � ��������� ���� ��������  ������, � ����������� �������������� ������ �� ����� ������  �� ����� ������ ����������� �������� ������� ����������� ��B�  ����� �������� �������.!�/B /Just L /Text ��������. ����   �������������� �����; ��������������.�������� ����������.�  ���������� ����� - �������� ��� ���������� �����; ��������  �������.�������� ����������.���������� ������������� - �� �  ����������� ���������� �������� ��� ���������� �������������   �������������, �������� ��� �����������; ��������������.��  ������� ����������.���������� ��������� - �������� ��� ����  ��������� ����������; ��������������.�������� �����.����� �  ����� - �������� ��� ����� �����; ��������������.���������   �����.����� ������������� - �� ����������� ���������� ����  ����� ��� ����� ������������ �������������, �������� ��� ���  ���������; ��������������.�������� �����.����� ��������� �  - �������� ��� ������������ �����. ����� ���� �������������  �� �������� �������� ��������� � ��� ������.!�� /B /Just L    /Text ����������� ���������� ��������. ��� ���� �� ������  ������ �����. ��������������.����������� ��� ���������� �6�  ����� ��������� ����������� ���������� - ���� ��� ���������  .��������. �������� � ���������� �������� � �����.!�k /B /  Just L /Text �������������� ����� ������������ ��������� ��  ���. ����������� ��� ����������� ����������.!��/B /Just L   /Text ��������� ��������� �����. �������� ��������� �����  � �������� ����� ������� ����, ��������� ������ ��������� �  ��������������, �������-���/�������� ������� �� ��������� �	  ���� ������� ���� ��� ������� ������� Control � ���������
  �� ���������. ��������������.��������.�� �������� ��� ��  ���; ��������������.��������.����������� ������������ - �  � ����������� ���������� �������� ������������ � ����������  � �������� ������; ��������������.��������.������������ ��  ���������� - �� ����������� ���������� �������� ����������  �� � ������������ �������� ������; ��������������.��������  .��������� - �������� ������������ �����-���� ���������� �  �������; ��������������.��������.��������� �������� - ����  ��. ��� ����� ������ ������ ���� �������� ����� ���� �����  ������� � ������� ������ ������. ���� �� ������ ��� ������,   �� ��� ������ �� ������ ��� �������� �� ������ ������� ���  ������ ����� ��������. ��� �����������  �� ��������� ������  ������ ��������� ���������������� �������� � ������ �������  ������ ���������� (������ �������� ������� ������, ������ -    �                                                            k. ��� ������ ��������� ��� ����� ������ ��������.��  
�   ������. ��������� ������ �� ��������� ����� � �������������  ����� k �����) �� ������ ����, ����� ���������� ������� ���   ���������). ��� ��������������� ��������� (�� n ���������       �  	  � 1050   �  ��Ab     �  �� L�   %  �  �  ������������� ����������� ������ [�     �  �� 	k#  v  -�   !�3 /T N /Just M /Text �������������� ����������� ��   ��!�% /H /Just L /Text �������� ��� �������!�� /B /Just L /  Text �������������� ������������ �������� � ������ ��������6  ���������� ����, ���������� ������ ���������. ��� ������ ��1   ������������ ��� �������� � �������������� ������ ��������$  �  ��� 
I - 4 M     � Topic@IDH_AssPCs  �    %  �  	  � 1051   �  ��;\     �  �� F�   "  � �������&  ��� ��������� ���������� U�     �  �� 	e~  �-�   !�0'   /T N /Just M /Text ���������� ��������� ��������!��/P /Ju(  st L /Text ��� ����� ���� ������� � ����� ���������� ������)  ��� ������������� �������� - �������� ������� "�������"  ��*  �������� ������ �������� �������. ������ � ������ ��������+     ������������� �� ���������� ������ ���������� ��������� ,  ��������. �������� ��������� �������� ����� ����������� ���-  � ������. ��� �������� ��� ������: "�������������", "�� ���.  ����������", "��������". ��� ����������� ������� ��������� /  ����� �������� ��������� �������. ��� ���� ���� ��� ��� ���0  �� ����������� ����������, �� ��� ����������� �� �����. ���!  �� ������� ���������� �������� ���� ��������, � ��������� �@  ����� ������ �����. ���������� ��������� �������� ���������A  �� ������ � ������� ������� (���������� �������� � ������ �2  ���� ������������� ��������� ����� ������������ ����� �����3  ������ �� ������ ������ ����� �������  . ��� ��������� ���    ����� ������� DEL, ���� ������ .  
� �                 5  . ������������ ���������� ����� ��� ���������� ������ � ���6   ������, ��� � ��� ��������.!�x /B /Just L /Text ��������7  ������� ������� ���� �� �������. ��� ���� ���������� ��� ��8  . ����������� �������   (������� ������ ���� ��������) ��� 9  ��.!�� /B /Just L /Text �������������� ���������� �������:  ��, � ������� ��������� ���������� ������������ � ���������;  �� ���������� ������, ����������� ��������� ��������� �����<  �� �������. ����������� �������   ��������� ������. ��� ��=  xt �������� ��� ���������!�� /B /Just L /Text �������� ���>   ����� ��������� ������ �������� �������.!�' /H /Just L /Te?  ��� ��������� ����������� ������ � ����. ��� ��������������P  ������). ����������� ������������� � ������ ������� �������C  �  ��� 
+ 1 8 Q     � Topic@IDH_CalcParams  �  D    �  	  � 1056   �  ��?`     �  �� J�   *  �% ���E  ������� ��������� ���������� ������� Y�     �  �� 	i� F   -�  
 !�8 /T N /Just M /Text ���������� ��������� ������Q  ���� �����!�� /P /Just L /Text ��������� ������ �������� ���  �	  �g�� 
: / 6 O     � Topic@IDH_Contents  �  �  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�        
� �                                                    I  ������ � �������������� � ���������� ����������� �����.��J  ������ ������������� ������������� �������������� ��� ���� K  ������� �, ���� ���� ������������� �������, �������������� L  .������� �������� ������ ������ ����� ����������� �� �����M  � ����, � �� ����� ������� ���������� ������������ ��������N  ������ � ������ ������� ������������ ����������� � �������O  � ������ ��� ���������� ��������� � �����.���� ������ ���� `  ����� ��������� ���� �������� ������ ��� ������� � ��������a  ���� ������������ ����� �� ����� � ������� ����������.!�/R  �� ����������� ���������� ���������� ��� ����� � ������� ��S  ������� �������.!�� /B /Just L /Text �������� ��� �����. T  ���� ����, ����� �������� ������� ������ ����� �������� ���U  ������.!�{ /B /Just L /Text ��������� �����������.  �����V  ���� ������. ������� ����� �������� ����� ������ �������� �W  ��� ����������� ������������� ��������� �� ����� ������ ���X  ��. ������ ������ �������� ���� ������� (1-2�), �� ��� ����Y  ������ ��� ������� ������������� ������������� ������������Z  �� � ������� ���� �������� � ������. ��  ������ ������� ��[   ����� ���������� ����� � �������. ��� ������ ������� �����\  � ���� ����������� ��������� �����, � �� ��������� ������ �]  � ��������������� �������������� ��� ��������� �������. ��^  ���.!�/B /Just L /Text ������ ������������� ������������_  ������� ����. � ������� ���� ����� ��������� ��������� ����p  B /Just L /Text �������� �����������. ��� ������������� �c  ��� �������� (����� � ����) ������������ �� ������ ����� (d  ������ ��������, ���� ����� ���� �������� �� ����� ������ ��  ��� �� ������ �� �������� ���� ��� �� ��� �������� ��������    ��������� ����� ������ �����.  
� �                     e  �� ����� ��������.!�C /B /Just L /Text ���������� �����. f  xt ��� �������� ��������. ��������� �� ����������� ��������g  ������ ��� �������������� �������� �����.!�[ /B /Just L /Teh  � ����������� ���������� ��������� ������������, ����������i  � ����� ����.!�� /B /Just L /Text ����������� ��������. �j  ���� ���������� ����� ���������������� ������������ �������k  �����. ����������� ���������� ����� � ��������, ������� ��l  ������ ��������������.!�� /B /Just L /Text �������� ����� m  ��� ������� ������ ��� ����������� �����, ��� ������� �����n  ���, ������������ ��� ������ � ������������ � ����������. o  ������ � ������������� ������ ���������� �� ����� ��������b  �-����� ����������;!�� /B /Just L /Text �� ����������� ����s  ���� ������ ����������� ������ �� ����������, ���� ����� �t  ��������� �� ����� ��� �� ����������, ���� � ������. ���� �u  ��������������� ����� ����� ����� ������������, �� ��������v  ��� �� �������� ����� � �������� .!�� /B /Just L /Text ���w  ���������� - ���� ��� ����� ����� ����� ������-������� ��x  �����-���. ����� ����� ��� ����� ����� ��������� ��������� y  ����� � �� ��� �� ��� ����� ��������� �� �����������.!�
 /Nz   /Just L!�G /I /Jump /Link f:\work\diplom\doc\adges.wmf /Ma{  cro /Play /Popup /Just C!�
 /N /Just L!�U /H /Just L /Text |  �� ��������� ����� ������������� ��������� ����������� � ��}  ��������:!�x /B /Just L /Text ����� ������ ���� �����������~   ������������ ����������� �� ����� � ������ �� �����-������  ����� � ������;!�^ /B /Just L /Text ��������� ����� ����� ��  ��������� ������ ����� � �� ������� ������ �� �������;!�O /q  B /Just L /Text ��������� ����������� ������ � ������� �����r   - ���� ����� ����� ������ ���������� � ����-����������. � �  ����� ������ ������ ������������� ����������� �����������, �  ���� ���������� �����������, ����������� ������ �������. ���  ���� ������ ����� ���������� ����� ���������� ����������� �  ��������������. �������� �� ����� ������������ �� �������� �  ����� � ��������. �������� ����-���������� ����� ���� ��� ��  �������� ������ � �������. ������ ����� ������������ �������  ��� ���� � ������ ����-���������� �� ���� ������� ����-�����  ������. ����� ����� ���� ������� � ����������. ������ ������   ������� �� ������ �����. ��������� ����� �������� ���������  � ���� ������� �� ���� � ������ ����-���������� � ���������  ��� ����-����� ���������� (�� �� ����-����������!). ������ �  ����-����� ���������� ��������� ����������� ������ ����� ��  ���. ����� ����-����� ����� �������� �������� � ����� ������  ������. ����������� �������� �� ����� ������������ ��� �����  �� � ����� � ����� ����:!�-/B /Just L /Text ������������  ����� �� ����� (����� ���� ����� ��������� ������ �����). �  ,  -\�� 
D 3 : S     � Topic@IDH_EditOfSchema  �    ������ �������� (��� � ����� �����).  
� �               �  ���� ������������� �������. ��������� ������ ������ ��������    ��� 
# . 5 N     � Topic@IDH_Schemes  �   �   �  	  � 3020   �  ��<]     �  �� G�     � ������  ������ ����� �������� V�     �  �� 	f  f-�   !�, /T�   N /Just M /Text ����������� ����� ������!� /H /Just L /T�  ext !�
 /N /Just L!�H /I /Jump /Link f:\work\diplom\doc\sch�  ema.wmf /Macro /Play /Popup /Just C!�
 /N /Just L!��/P /Ju�  st L /Text �����  ������� �� ����� ���� ����� (��������� � �  ����� ����������) � ������. �������� ������ ����������� ���  ��� ���� ��������� ������� ����������, ���������������� ����   ��������� ������������ ���������� ������� ����. �����-�����  ������� ������������� ���� � �����. ��������� ������ �������  ������ � ������� �� ����� � ������, � ������ ������������� �   /Text ������������������ �������� ����� �������� ����� ���  Just L /Text ��� ���� ������������ ��������� ���������� ����  �� ������������ ��������� ������������ �����������;!�J /B /�  , ������������� ���������������;!�J /B /Just L /Text ��� ���  �� �������:!�K /B /Just L /Text ��� ������������� ���������  �� ������-������������. ����������� ������ ����������� � ��  ��� ������� ������ ���������������� ����-���������� � ������  �����, ���������������� ������������) ����������� �� �������  ������ � ���� ������ (������������, ���������������� ������  �� ��������������� ����������� ������������� ��� ������. ��  �������������� ����������� � ������� ������ � �������������  ������� �������������� ���� �����. �������� ������� �� �����  ���� ����������� ����� � ������ �������������� � ����������  	  � 1057   �  ��7X     �  �� B�   "  � ������ �����  �� ����������������� Q�     �  �� 	a�  �-�   !�0 /T �  N /Just M /Text ������ ������ ���������������!�)/P /Just L�  ����������.!��/P /Just L /Text ��� ������������� � ������    ���� ��������� ������� ������� � ������.  
� �           �  ���������, ������� �������������, � ������ ������ ������ ��  ����� �������. � ��������� ������, ���� ��� �������������� �  ������������ � � ���������� �� ���� ���������� ���� ��������   ������������ ��������� �������������� ����� ��������, ��� �  �� ����� ����������� �������� �������� ���������������. ����  ������� ���������-��. ����� ��������� � ������ ������������  � ������������� ������ �� ������������� ����� � ��� ��������  ���������� � ������������ ������ � �������, � �������� �����  � � ������ �������� ����� � ������ ����-����������. ������ �  �������� ������. ���������������� �� ������ ���� ����������  ��������������� ���������� �������) ����������� � ����� ���  ��������� ������ (��� ������������� �������� �� ������, �� �  � (���������� ��������������� � �������������� ���������). �  ������� ������� ����� ����������� ���������-������ ��������6�  �  ��� 
F ) 0 I     � Topic@IDH_PE  �    �                                                                 �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                             �                                                                 !�  !�  !�  !�                                             �  �  �N�� 
G 0 7 P     � Topic@IDH_Interface  �  